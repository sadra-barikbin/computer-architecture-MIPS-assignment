library verilog;
use verilog.vl_types.all;
entity Instruction_memory is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        address         : in     vl_logic_vector(31 downto 0);
        data_out        : out    vl_logic_vector(31 downto 0)
    );
end Instruction_memory;
