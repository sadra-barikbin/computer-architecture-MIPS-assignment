library verilog;
use verilog.vl_types.all;
entity self_test is
end self_test;
