library verilog;
use verilog.vl_types.all;
entity mips_tester is
end mips_tester;
