library verilog;
use verilog.vl_types.all;
entity MIPS is
    port(
        CLOCK_27        : in     vl_logic;
        CLOCK_50        : in     vl_logic;
        EXT_CLOCK       : in     vl_logic;
        KEY             : in     vl_logic_vector(3 downto 0);
        SW              : in     vl_logic_vector(17 downto 0);
        HEX0            : out    vl_logic_vector(6 downto 0);
        HEX1            : out    vl_logic_vector(6 downto 0);
        HEX2            : out    vl_logic_vector(6 downto 0);
        HEX3            : out    vl_logic_vector(6 downto 0);
        HEX4            : out    vl_logic_vector(6 downto 0);
        HEX5            : out    vl_logic_vector(6 downto 0);
        HEX6            : out    vl_logic_vector(6 downto 0);
        HEX7            : out    vl_logic_vector(6 downto 0);
        LEDG            : out    vl_logic_vector(8 downto 0);
        LEDR            : out    vl_logic_vector(17 downto 0);
        DRAM_DQ         : inout  vl_logic_vector(15 downto 0);
        DRAM_ADDR       : out    vl_logic_vector(11 downto 0);
        DRAM_LDQM       : out    vl_logic;
        DRAM_UDQM       : out    vl_logic;
        DRAM_WE_N       : out    vl_logic;
        DRAM_CAS_N      : out    vl_logic;
        DRAM_RAS_N      : out    vl_logic;
        DRAM_CS_N       : out    vl_logic;
        DRAM_BA_0       : out    vl_logic;
        DRAM_BA_1       : out    vl_logic;
        DRAM_CLK        : out    vl_logic;
        DRAM_CKE        : out    vl_logic;
        FL_DQ           : inout  vl_logic_vector(7 downto 0);
        FL_ADDR         : out    vl_logic_vector(21 downto 0);
        FL_WE_N         : out    vl_logic;
        FL_RST_N        : out    vl_logic;
        FL_OE_N         : out    vl_logic;
        FL_CE_N         : out    vl_logic;
        SRAM_DQ         : inout  vl_logic_vector(15 downto 0);
        SRAM_ADDR       : out    vl_logic_vector(17 downto 0);
        SRAM_UB_N       : out    vl_logic;
        SRAM_LB_N       : out    vl_logic;
        SRAM_WE_N       : out    vl_logic;
        SRAM_CE_N       : out    vl_logic;
        SRAM_OE_N       : out    vl_logic;
        OTG_DATA        : inout  vl_logic_vector(15 downto 0);
        OTG_ADDR        : out    vl_logic_vector(1 downto 0);
        OTG_CS_N        : out    vl_logic;
        OTG_RD_N        : out    vl_logic;
        OTG_WR_N        : out    vl_logic;
        OTG_RST_N       : out    vl_logic;
        OTG_FSPEED      : out    vl_logic;
        OTG_LSPEED      : out    vl_logic;
        OTG_INT0        : in     vl_logic;
        OTG_INT1        : in     vl_logic;
        OTG_DREQ0       : in     vl_logic;
        OTG_DREQ1       : in     vl_logic;
        OTG_DACK0_N     : out    vl_logic;
        OTG_DACK1_N     : out    vl_logic;
        LCD_ON          : out    vl_logic;
        LCD_BLON        : out    vl_logic;
        LCD_RW          : out    vl_logic;
        LCD_EN          : out    vl_logic;
        LCD_RS          : out    vl_logic;
        LCD_DATA        : inout  vl_logic_vector(7 downto 0);
        TDI             : in     vl_logic;
        TCK             : in     vl_logic;
        TCS             : in     vl_logic;
        TDO             : out    vl_logic;
        I2C_SDAT        : inout  vl_logic;
        I2C_SCLK        : out    vl_logic;
        PS2_DAT         : in     vl_logic;
        PS2_CLK         : in     vl_logic;
        VGA_CLK         : out    vl_logic;
        VGA_HS          : out    vl_logic;
        VGA_VS          : out    vl_logic;
        VGA_BLANK       : out    vl_logic;
        VGA_SYNC        : out    vl_logic;
        VGA_R           : out    vl_logic_vector(9 downto 0);
        VGA_G           : out    vl_logic_vector(9 downto 0);
        VGA_B           : out    vl_logic_vector(9 downto 0);
        ENET_DATA       : inout  vl_logic_vector(15 downto 0);
        ENET_CMD        : out    vl_logic;
        ENET_CS_N       : out    vl_logic;
        ENET_WR_N       : out    vl_logic;
        ENET_RD_N       : out    vl_logic;
        ENET_RST_N      : out    vl_logic;
        ENET_INT        : in     vl_logic;
        ENET_CLK        : out    vl_logic;
        AUD_ADCLRCK     : inout  vl_logic;
        AUD_ADCDAT      : in     vl_logic;
        AUD_DACLRCK     : inout  vl_logic;
        AUD_DACDAT      : out    vl_logic;
        AUD_BCLK        : inout  vl_logic;
        AUD_XCK         : out    vl_logic;
        TD_DATA         : in     vl_logic_vector(7 downto 0);
        TD_HS           : in     vl_logic;
        TD_VS           : in     vl_logic;
        TD_RESET        : out    vl_logic;
        TD_CLK27        : in     vl_logic;
        GPIO_0          : inout  vl_logic_vector(35 downto 0);
        GPIO_1          : inout  vl_logic_vector(35 downto 0)
    );
end MIPS;
